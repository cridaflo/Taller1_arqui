module MI_ROM #(parameter DATA_BUS_IN = 11, parameter DATA_BUS_OUT = 44)(BUS_IN, BUS_OUT,CLK);

//=======================================================
//  PORT declarations
//=======================================================
output BUS_OUT [DATA_BUS_OUT-1: 0];
input BUS_IN [DATA_BUS_IN-1:0];
input CLK;
//=======================================================
//  Structural coding
//=======================================================


// REGISTER : SEQUENTIAL
	always @ ( negedge CLK) begin
		case (Bus_IN)
		//inicializa
			4'd0000:BUS_OUT <= 41'b10000010000000101010010100000000000000;
			4'd0001:BUS_OUT <= 41'b00000000000000000000010111100000000000;
		//addcc
			4'd1600:BUS_OUT <= 41'b00000000000000000000010110111001000010;
			4'd1601:BUS_OUT <= 41'b00000100000100000100001111011111111111;
			4'd1602:BUS_OUT <= 41'b10101000000000001000110000000000000000;
			4'd1603:BUS_OUT <= 41'b00000110001000000100001111011111111111;
		//arncc
			4'd1624:BUS_OUT <= 41'b00000000000000000000010110111001011010;
			4'd1625:BUS_OUT <= 41'b00000100000100000100001011011111111111;
			4'd1626:BUS_OUT <= 41'b10101000000000001000101100000000000000;
			4'd1627:BUS_OUT <= 41'b00000110001000000100001011011111111111;

		//branching
			4'd0002:BUS_OUT <= 41'b10101000000010001000101000000000000000;
			4'd0003:BUS_OUT <= 41'b10001000000010001000111100000000000000;
			4'd0004:BUS_OUT <= 41'b10001000000010001000111100000000000000;
			4'd0005:BUS_OUT <= 41'b10101000000010101000111100000000000000;
			4'd0006:BUS_OUT <= 41'b10101000000010101000111100000000000000;
			4'd0007:BUS_OUT <= 41'b10101000000010101000111100000000000000;
			4'd0008:BUS_OUT <= 41'b10101010100010101000100010100000001100;
			4'd0009:BUS_OUT <= 41'b10101010100010101000100010100000001101;
			4'd0010:BUS_OUT <= 41'b10101010100010101000100001000000001100;
			4'd0011:BUS_OUT <= 41'b00000000000000000000010111011111111111;
			4'd0012:BUS_OUT <= 41'b10000010001010000000100011000000000000;
			4'd0013:BUS_OUT <= 41'b10101010101010101000100010100000010000;
			4'd0014:BUS_OUT <= 41'b00000000000000000000010110000000001100;
			4'd0015:BUS_OUT <= 41'b00000000000000000000010111011111111111;
			4'd0016:BUS_OUT <= 41'b00000000000000000000010110100000010011;
			4'd0017:BUS_OUT <= 41'b00000000000000000000010100100000001100;
			4'd0018:BUS_OUT <= 41'b00000000000000000000010111011111111111;
			4'd0019:BUS_OUT <= 41'b00000000000000000000010101100000001100;
			4'd0020:BUS_OUT <= 41'b00000000000000000000010111011111111111:
			
		//incremntar pc
		   4'd2047:BUS_OUT <= 41'b10000000000010000000111011000000000000;
			
			
		endcase
	end;