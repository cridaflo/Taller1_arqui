module programMem #(parameter DATAWIDTH_BUS=32)(
// ------------- Inputs ---------------
   BusDirecciones,
 
// ------------ Outputs ---------------
 
	BusDatos
);
 
//=======================================================
//  PARAMETER declarations
//=======================================================
 
 
//=======================================================
//  PORT declarations
//=======================================================
input [DATAWIDTH_BUS-1:0] BusDirecciones; 
output reg [DATAWIDTH_BUS-1:0] BusDatos; 
 
 
//=======================================================
//  REG/WIRE declarations
//=======================================================
 
 
 
//=======================================================
//  Structural coding
//=======================================================
 always @(*)
 begin
	case (BusDirecciones)
	32'b0000000000000000000100000000000: BusDatos=32'b10000010100000000010000000000001;
	32'b0000000000000000000100000000001: BusDatos=32'b10000100100000000010000000000001;
	32'b0000000000000000000100000000010: BusDatos=32'b10000110100000000010000000000000;
	32'b0000000000000000000100000000011: BusDatos=32'b10001000100000000011111111110110;
	32'b0000000000000000000100000000100: BusDatos=32'b10000010100000001000000000000011;
	32'b0000000000000000000100000000101: BusDatos=32'b10000110100000001000000000000000;
	32'b0000000000000000000100000000110: BusDatos=32'b10000100100000000100000000000000;
	32'b0000000000000000000100000000111: BusDatos=32'b00001100101111111111111111111100;
	32'b0000000000000000000100000001000: BusDatos=32'b10000010100000001110000000000000;
	32'b0000000000000000000100000001001: BusDatos=32'b10000110101100001100000000000011;
	32'b0000000000000000000100000001010: BusDatos=32'b10000110100000001100000000000010;
	32'b0000000000000000000100000001011: BusDatos=32'b00000010100000000000000000000011;
	32'b0000000000000000000100000001100: BusDatos=32'b10000100100000000110000000000000;
	32'b0000000000000000000100000001101: BusDatos=32'b00010000101111111111111111111011;
	32'b0000000000000000000100000001110: BusDatos=32'b00000000000000000000000000000000;
	default: BusDatos=32'b00000000000000000000000000000000;
	endcase
	end
 
endmodule
