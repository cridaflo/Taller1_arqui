//=======================================================
//  MODULE Definition
//=======================================================
module CC_MUX_REG #(parameter DATAWIDTH_DECODER_OUT=38, parameter DATAWIDTH_BUS=32)(
	//////////// OUTPUTS //////////
	CC_MUX_REG_TO_BUS_OUT,
	//////////// INPUTS //////////
	CC_MUX_REG_R0,
	CC_MUX_REG_R1,
	CC_MUX_REG_R2,
	CC_MUX_REG_R3,
	CC_MUX_REG_R4,
	CC_MUX_REG_R5,
	CC_MUX_REG_R6,
	CC_MUX_REG_R7,
	CC_MUX_REG_R8,
	CC_MUX_REG_R9,
	CC_MUX_REG_R10,
	CC_MUX_REG_R11,
	CC_MUX_REG_R12,
	CC_MUX_REG_R13,
	CC_MUX_REG_R14,
	CC_MUX_REG_R15,
	CC_MUX_REG_R16,
	CC_MUX_REG_R17,
	CC_MUX_REG_R18,
	CC_MUX_REG_R19,
	CC_MUX_REG_R20,
	CC_MUX_REG_R21,
	CC_MUX_REG_R22,
	CC_MUX_REG_R23,
	CC_MUX_REG_R24,
	CC_MUX_REG_R25,
	CC_MUX_REG_R26,
	CC_MUX_REG_R27,
	CC_MUX_REG_R28,
	CC_MUX_REG_R29,
	CC_MUX_REG_R30,
	CC_MUX_REG_R31,
	CC_MUX_REG_R32,
	CC_MUX_REG_R33,
	CC_MUX_REG_R34,
	CC_MUX_REG_R35,
	CC_MUX_REG_R36,
	CC_MUX_REG_R37,
	CC_MUX_REG_DECOD_SELECTION
);
//=======================================================
//  PARAMETER declarations
//=======================================================

//=======================================================
//  PORT declarations
//=======================================================
   output reg [DATAWIDTH_BUS-1:0]CC_MUX_REG_TO_BUS_OUT;
	input [DATAWIDTH_BUS-1:0]CC_MUX_REG_R0;
	input [DATAWIDTH_BUS-1:0]CC_MUX_REG_R1;
	input [DATAWIDTH_BUS-1:0]CC_MUX_REG_R2;
	input [DATAWIDTH_BUS-1:0]CC_MUX_REG_R3;
	input [DATAWIDTH_BUS-1:0]CC_MUX_REG_R4;
	input [DATAWIDTH_BUS-1:0]CC_MUX_REG_R5;
	input [DATAWIDTH_BUS-1:0]CC_MUX_REG_R6;
	input [DATAWIDTH_BUS-1:0]CC_MUX_REG_R7;
	input [DATAWIDTH_BUS-1:0]CC_MUX_REG_R8;
	input [DATAWIDTH_BUS-1:0]CC_MUX_REG_R9;
	input [DATAWIDTH_BUS-1:0]CC_MUX_REG_R10;
	input [DATAWIDTH_BUS-1:0]CC_MUX_REG_R11;
	input [DATAWIDTH_BUS-1:0]CC_MUX_REG_R12;
	input [DATAWIDTH_BUS-1:0]CC_MUX_REG_R13;
	input [DATAWIDTH_BUS-1:0]CC_MUX_REG_R14;
	input [DATAWIDTH_BUS-1:0]CC_MUX_REG_R15;
	input [DATAWIDTH_BUS-1:0]CC_MUX_REG_R16;
	input [DATAWIDTH_BUS-1:0]CC_MUX_REG_R17;
	input [DATAWIDTH_BUS-1:0]CC_MUX_REG_R18;
	input [DATAWIDTH_BUS-1:0]CC_MUX_REG_R19;
	input [DATAWIDTH_BUS-1:0]CC_MUX_REG_R20;
	input [DATAWIDTH_BUS-1:0]CC_MUX_REG_R21;
	input [DATAWIDTH_BUS-1:0]CC_MUX_REG_R22;
	input [DATAWIDTH_BUS-1:0]CC_MUX_REG_R23;
	input [DATAWIDTH_BUS-1:0]CC_MUX_REG_R24;
	input [DATAWIDTH_BUS-1:0]CC_MUX_REG_R25;
	input [DATAWIDTH_BUS-1:0]CC_MUX_REG_R26;
	input [DATAWIDTH_BUS-1:0]CC_MUX_REG_R27;
	input [DATAWIDTH_BUS-1:0]CC_MUX_REG_R28;
	input [DATAWIDTH_BUS-1:0]CC_MUX_REG_R29;
	input [DATAWIDTH_BUS-1:0]CC_MUX_REG_R30;
	input [DATAWIDTH_BUS-1:0]CC_MUX_REG_R31;
	input [DATAWIDTH_BUS-1:0]CC_MUX_REG_R32;
	input [DATAWIDTH_BUS-1:0]CC_MUX_REG_R33;
	input [DATAWIDTH_BUS-1:0]CC_MUX_REG_R34;
	input [DATAWIDTH_BUS-1:0]CC_MUX_REG_R35;
	input [DATAWIDTH_BUS-1:0]CC_MUX_REG_R36;
	input [DATAWIDTH_BUS-1:0]CC_MUX_REG_R37;
	input [DATAWIDTH_DECODER_OUT-1:0]CC_MUX_REG_DECOD_SELECTION;
//=======================================================
//  REG/WIRE declarations
//=======================================================

//=======================================================
//  Structural coding
//=======================================================
//INPUT LOGIC: COMBINATIONAL
	always@(*)
	begin
	case (CC_MUX_REG_DECOD_SELECTION)
		38'b00000000000000000000000000000000000001: CC_MUX_REG_TO_BUS_OUT = CC_MUX_REG_R0;
		38'b00000000000000000000000000000000000010: CC_MUX_REG_TO_BUS_OUT = CC_MUX_REG_R1;
		38'b00000000000000000000000000000000000100: CC_MUX_REG_TO_BUS_OUT = CC_MUX_REG_R2;
		38'b00000000000000000000000000000000001000: CC_MUX_REG_TO_BUS_OUT = CC_MUX_REG_R3;
		38'b00000000000000000000000000000000010000: CC_MUX_REG_TO_BUS_OUT = CC_MUX_REG_R4;
		38'b00000000000000000000000000000000100000: CC_MUX_REG_TO_BUS_OUT = CC_MUX_REG_R5;
		38'b00000000000000000000000000000001000000: CC_MUX_REG_TO_BUS_OUT = CC_MUX_REG_R6;
		38'b00000000000000000000000000000010000000: CC_MUX_REG_TO_BUS_OUT = CC_MUX_REG_R7;
		38'b00000000000000000000000000000100000000: CC_MUX_REG_TO_BUS_OUT = CC_MUX_REG_R8;
		38'b00000000000000000000000000001000000000: CC_MUX_REG_TO_BUS_OUT = CC_MUX_REG_R9;
		38'b00000000000000000000000000010000000000: CC_MUX_REG_TO_BUS_OUT = CC_MUX_REG_R10;
		38'b00000000000000000000000000100000000000: CC_MUX_REG_TO_BUS_OUT = CC_MUX_REG_R11;
		38'b00000000000000000000000001000000000000: CC_MUX_REG_TO_BUS_OUT = CC_MUX_REG_R12;
		38'b00000000000000000000000010000000000000: CC_MUX_REG_TO_BUS_OUT = CC_MUX_REG_R13;
		38'b00000000000000000000000100000000000000: CC_MUX_REG_TO_BUS_OUT = CC_MUX_REG_R14;
		38'b00000000000000000000001000000000000000: CC_MUX_REG_TO_BUS_OUT = CC_MUX_REG_R15;
		38'b00000000000000000000010000000000000000: CC_MUX_REG_TO_BUS_OUT = CC_MUX_REG_R16;
		38'b00000000000000000000100000000000000000: CC_MUX_REG_TO_BUS_OUT = CC_MUX_REG_R17;
		38'b00000000000000000001000000000000000000: CC_MUX_REG_TO_BUS_OUT = CC_MUX_REG_R18;
		38'b00000000000000000010000000000000000000: CC_MUX_REG_TO_BUS_OUT = CC_MUX_REG_R19;
		38'b00000000000000000100000000000000000000: CC_MUX_REG_TO_BUS_OUT = CC_MUX_REG_R20;
		38'b00000000000000001000000000000000000000: CC_MUX_REG_TO_BUS_OUT = CC_MUX_REG_R21;
		38'b00000000000000010000000000000000000000: CC_MUX_REG_TO_BUS_OUT = CC_MUX_REG_R22;
		38'b00000000000000100000000000000000000000: CC_MUX_REG_TO_BUS_OUT = CC_MUX_REG_R23;
		38'b00000000000001000000000000000000000000: CC_MUX_REG_TO_BUS_OUT = CC_MUX_REG_R24;
		38'b00000000000010000000000000000000000000: CC_MUX_REG_TO_BUS_OUT = CC_MUX_REG_R25;
		38'b00000000000100000000000000000000000000: CC_MUX_REG_TO_BUS_OUT = CC_MUX_REG_R26;
		38'b00000000001000000000000000000000000000: CC_MUX_REG_TO_BUS_OUT = CC_MUX_REG_R27;
		38'b00000000010000000000000000000000000000: CC_MUX_REG_TO_BUS_OUT = CC_MUX_REG_R28;
		38'b00000000100000000000000000000000000000: CC_MUX_REG_TO_BUS_OUT = CC_MUX_REG_R29;
		38'b00000001000000000000000000000000000000: CC_MUX_REG_TO_BUS_OUT = CC_MUX_REG_R30;
		38'b00000010000000000000000000000000000000: CC_MUX_REG_TO_BUS_OUT = CC_MUX_REG_R31;
		38'b00000100000000000000000000000000000000: CC_MUX_REG_TO_BUS_OUT = CC_MUX_REG_R32;
		38'b00001000000000000000000000000000000000: CC_MUX_REG_TO_BUS_OUT = CC_MUX_REG_R33;
		38'b00010000000000000000000000000000000000: CC_MUX_REG_TO_BUS_OUT = CC_MUX_REG_R34;
		38'b00100000000000000000000000000000000000: CC_MUX_REG_TO_BUS_OUT = CC_MUX_REG_R35;
		38'b01000000000000000000000000000000000000: CC_MUX_REG_TO_BUS_OUT = CC_MUX_REG_R36;
		38'b10000000000000000000000000000000000000: CC_MUX_REG_TO_BUS_OUT = CC_MUX_REG_R37;
		default : CC_MUX_REG_TO_BUS_OUT = 0;
		endcase
	end
endmodule
