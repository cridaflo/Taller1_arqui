module programMem #(parameter DATAWIDTH_BUS = 32)(
// ------------- Inputs ---------------
   RD,
	WR,
	BusDirecciones,
 
// ------------ Outputs ---------------
 
	BusDatos
);
 
//=======================================================
//  PARAMETER declarations
//=======================================================
 
 
//=======================================================
//  PORT declarations
//=======================================================
input RD;
input WR;
input [DATAWIDTH_BUS-1:0] BusDirecciones; 
output reg [DATAWIDTH_BUS-1:0] BusDatos; 
 
 
//=======================================================
//  REG/WIRE declarations
//=======================================================
 
reg [DATAWIDTH_BUS-1:0] BusMemoria;
 
//=======================================================
//  Structural coding
//=======================================================
 always @(*)
 begin
 if (RD==0)
		BusMemoria <= 32'b00000000000000000000000000000000;
	else
		BusMemoria <= BusDirecciones; 
	case (BusMemoria)
	32'b0000000000000000000100000000000: BusDatos=32'b10000010100000000010000000000001; //addcc %r0, 1, %r1   
	32'b0000000000000000000100000000100: BusDatos=32'b10000100100000000010000000000001; //addcc %r0, 1, %r2 
	32'b0000000000000000000100000001000: BusDatos=32'b10000110100000000010000000000000; //addcc %r0, 0, %r3 
	32'b0000000000000000000100000001100: BusDatos=32'b10001000100000000011111111110110; //addcc %r0, -10, %r4 
	32'b0000000000000000000100000010000: BusDatos=32'b10000010100000001000000000000011; //addcc %r2, %r3, %r1
	32'b0000000000000000000100000010100: BusDatos=32'b10000110100000001000000000000000; //addcc %r2, %r0, %r3
	32'b0000000000000000000100000011000: BusDatos=32'b10000100100000000100000000000000; //addcc %r1, %r0, %r2
	32'b0000000000000000000100000011100: BusDatos=32'b10001000100000010010000000000001; //addcc %r4, 1, %r4 
	32'b0000000000000000000100000100000: BusDatos=32'b00001100101111111111111111110000; //bneg -4 		
	32'b0000000000000000000100000100100: BusDatos=32'b10000010100000001110000000000000; //addcc %r3, 0, %r1 
	32'b0000000000000000000100000101000: BusDatos=32'b10000110101100001100000000000011; //orncc %r3, %r3, %r3 
	32'b0000000000000000000100000101100: BusDatos=32'b10000110100000001110000000000001; //adcc %r3, 1, %r3
	32'b0000000000000000000100000110000: BusDatos=32'b10000110100000001100000000000010; //addcc %r3, %r2, %r3
	32'b0000000000000000000100000110100: BusDatos=32'b00000010100000000000000000001100; //be 3 
	32'b0000000000000000000100000111000: BusDatos=32'b10000100100000000110000000000000; //addcc %r1, 0, %r2
	32'b0000000000000000000100000111100: BusDatos=32'b00010000101111111111111111101000; // ba -6
        32'b0000000000000000000100001000000: BusDatos=32'b00000000000000000000000000000000; //fin
	default: BusDatos=32'b00000000000000000000000000000000;
	endcase
end
endmodule
