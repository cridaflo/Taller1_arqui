//=======================================================
//  MODULE Definition
//=======================================================
module CC_MUX_REG #(parameter DATAWIDTH_DECODER_OUT=38, parameter DATAWIDTH_BUS=32)(
	//////////// OUTPUTS //////////
	CC_MUX_REG_TO_BUS_OUT,
	//////////// INPUTS //////////
	REG_TO_MUX_R0,
	REG_TO_MUX_R1,
	REG_TO_MUX_R2,
	REG_TO_MUX_R3,
	REG_TO_MUX_R4,
	REG_TO_MUX_R5,
	REG_TO_MUX_R6,
	REG_TO_MUX_R7,
	REG_TO_MUX_R8,
	REG_TO_MUX_R9,
	REG_TO_MUX_R10,
	REG_TO_MUX_R11,
	REG_TO_MUX_R12,
	REG_TO_MUX_R13,
	REG_TO_MUX_R14,
	REG_TO_MUX_R15,
	REG_TO_MUX_R16,
	REG_TO_MUX_R17,
	REG_TO_MUX_R18,
	REG_TO_MUX_R19,
	REG_TO_MUX_R20,
	REG_TO_MUX_R21,
	REG_TO_MUX_R22,
	REG_TO_MUX_R23,
	REG_TO_MUX_R24,
	REG_TO_MUX_R25,
	REG_TO_MUX_R26,
	REG_TO_MUX_R27,
	REG_TO_MUX_R28,
	REG_TO_MUX_R29,
	REG_TO_MUX_R30,
	REG_TO_MUX_R31,
	REG_TO_MUX_R32,
	REG_TO_MUX_R33,
	REG_TO_MUX_R34,
	REG_TO_MUX_R35,
	REG_TO_MUX_R36,
	REG_TO_MUX_R37,
	CC_MUX_REG_DECOD_SELECTION
);
//=======================================================
//  PARAMETER declarations
//=======================================================

//=======================================================
//  PORT declarations
//=======================================================
   output reg [DATAWIDTH_BUS-1:0]CC_MUX_REG_TO_BUS_OUT;
	input [DATAWIDTH_BUS-1:0]REG_TO_MUX_R0;
	input [DATAWIDTH_BUS-1:0]REG_TO_MUX_R1;
	input [DATAWIDTH_BUS-1:0]REG_TO_MUX_R2;
	input [DATAWIDTH_BUS-1:0]REG_TO_MUX_R3;
	input [DATAWIDTH_BUS-1:0]REG_TO_MUX_R4;
	input [DATAWIDTH_BUS-1:0]REG_TO_MUX_R5;
	input [DATAWIDTH_BUS-1:0]REG_TO_MUX_R6;
	input [DATAWIDTH_BUS-1:0]REG_TO_MUX_R7;
	input [DATAWIDTH_BUS-1:0]REG_TO_MUX_R8;
	input [DATAWIDTH_BUS-1:0]REG_TO_MUX_R9;
	input [DATAWIDTH_BUS-1:0]REG_TO_MUX_R10;
	input [DATAWIDTH_BUS-1:0]REG_TO_MUX_R11;
	input [DATAWIDTH_BUS-1:0]REG_TO_MUX_R12;
	input [DATAWIDTH_BUS-1:0]REG_TO_MUX_R13;
	input [DATAWIDTH_BUS-1:0]REG_TO_MUX_R14;
	input [DATAWIDTH_BUS-1:0]REG_TO_MUX_R15;
	input [DATAWIDTH_BUS-1:0]REG_TO_MUX_R16;
	input [DATAWIDTH_BUS-1:0]REG_TO_MUX_R17;
	input [DATAWIDTH_BUS-1:0]REG_TO_MUX_R18;
	input [DATAWIDTH_BUS-1:0]REG_TO_MUX_R19;
	input [DATAWIDTH_BUS-1:0]REG_TO_MUX_R20;
	input [DATAWIDTH_BUS-1:0]REG_TO_MUX_R21;
	input [DATAWIDTH_BUS-1:0]REG_TO_MUX_R22;
	input [DATAWIDTH_BUS-1:0]REG_TO_MUX_R23;
	input [DATAWIDTH_BUS-1:0]REG_TO_MUX_R24;
	input [DATAWIDTH_BUS-1:0]REG_TO_MUX_R25;
	input [DATAWIDTH_BUS-1:0]REG_TO_MUX_R26;
	input [DATAWIDTH_BUS-1:0]REG_TO_MUX_R27;
	input [DATAWIDTH_BUS-1:0]REG_TO_MUX_R28;
	input [DATAWIDTH_BUS-1:0]REG_TO_MUX_R29;
	input [DATAWIDTH_BUS-1:0]REG_TO_MUX_R30;
	input [DATAWIDTH_BUS-1:0]REG_TO_MUX_R31;
	input [DATAWIDTH_BUS-1:0]REG_TO_MUX_R32;
	input [DATAWIDTH_BUS-1:0]REG_TO_MUX_R33;
	input [DATAWIDTH_BUS-1:0]REG_TO_MUX_R34;
	input [DATAWIDTH_BUS-1:0]REG_TO_MUX_R35;
	input [DATAWIDTH_BUS-1:0]REG_TO_MUX_R36;
	input [DATAWIDTH_BUS-1:0]REG_TO_MUX_R37;
	input [DATAWIDTH_DECODER_OUT-1:0]CC_MUX_REG_DECOD_SELECTION;
//=======================================================
//  REG/WIRE declarations
//=======================================================

//=======================================================
//  Structural coding
//=======================================================
//INPUT LOGIC: COMBINATIONAL
	always@(*)
	begin
	case (CC_MUX_REG_DECOD_SELECTION)
		38'b00000000000000000000000000000000000001: CC_MUX_REG_TO_BUS_OUT = REG_TO_MUX_R0;
		38'b00000000000000000000000000000000000010: CC_MUX_REG_TO_BUS_OUT = REG_TO_MUX_R1;
		38'b00000000000000000000000000000000000100: CC_MUX_REG_TO_BUS_OUT = REG_TO_MUX_R2;
		38'b00000000000000000000000000000000001000: CC_MUX_REG_TO_BUS_OUT = REG_TO_MUX_R3;
		38'b00000000000000000000000000000000010000: CC_MUX_REG_TO_BUS_OUT = REG_TO_MUX_R4;
		38'b00000000000000000000000000000000100000: CC_MUX_REG_TO_BUS_OUT = REG_TO_MUX_R5;
		38'b00000000000000000000000000000001000000: CC_MUX_REG_TO_BUS_OUT = REG_TO_MUX_R6;
		38'b00000000000000000000000000000010000000: CC_MUX_REG_TO_BUS_OUT = REG_TO_MUX_R7;
		38'b00000000000000000000000000000100000000: CC_MUX_REG_TO_BUS_OUT = REG_TO_MUX_R8;
		38'b00000000000000000000000000001000000000: CC_MUX_REG_TO_BUS_OUT = REG_TO_MUX_R9;
		38'b00000000000000000000000000010000000000: CC_MUX_REG_TO_BUS_OUT = REG_TO_MUX_R10;
		38'b00000000000000000000000000100000000000: CC_MUX_REG_TO_BUS_OUT = REG_TO_MUX_R11;
		38'b00000000000000000000000001000000000000: CC_MUX_REG_TO_BUS_OUT = REG_TO_MUX_R12;
		38'b00000000000000000000000010000000000000: CC_MUX_REG_TO_BUS_OUT = REG_TO_MUX_R13;
		38'b00000000000000000000000100000000000000: CC_MUX_REG_TO_BUS_OUT = REG_TO_MUX_R14;
		38'b00000000000000000000001000000000000000: CC_MUX_REG_TO_BUS_OUT = REG_TO_MUX_R15;
		38'b00000000000000000000010000000000000000: CC_MUX_REG_TO_BUS_OUT = REG_TO_MUX_R16;
		38'b00000000000000000000100000000000000000: CC_MUX_REG_TO_BUS_OUT = REG_TO_MUX_R17;
		38'b00000000000000000001000000000000000000: CC_MUX_REG_TO_BUS_OUT = REG_TO_MUX_R18;
		38'b00000000000000000010000000000000000000: CC_MUX_REG_TO_BUS_OUT = REG_TO_MUX_R19;
		38'b00000000000000000100000000000000000000: CC_MUX_REG_TO_BUS_OUT = REG_TO_MUX_R20;
		38'b00000000000000001000000000000000000000: CC_MUX_REG_TO_BUS_OUT = REG_TO_MUX_R21;
		38'b00000000000000010000000000000000000000: CC_MUX_REG_TO_BUS_OUT = REG_TO_MUX_R22;
		38'b00000000000000100000000000000000000000: CC_MUX_REG_TO_BUS_OUT = REG_TO_MUX_R23;
		38'b00000000000001000000000000000000000000: CC_MUX_REG_TO_BUS_OUT = REG_TO_MUX_R24;
		38'b00000000000010000000000000000000000000: CC_MUX_REG_TO_BUS_OUT = REG_TO_MUX_R25;
		38'b00000000000100000000000000000000000000: CC_MUX_REG_TO_BUS_OUT = REG_TO_MUX_R26;
		38'b00000000001000000000000000000000000000: CC_MUX_REG_TO_BUS_OUT = REG_TO_MUX_R27;
		38'b00000000010000000000000000000000000000: CC_MUX_REG_TO_BUS_OUT = REG_TO_MUX_R28;
		38'b00000000100000000000000000000000000000: CC_MUX_REG_TO_BUS_OUT = REG_TO_MUX_R29;
		38'b00000001000000000000000000000000000000: CC_MUX_REG_TO_BUS_OUT = REG_TO_MUX_R30;
		38'b00000010000000000000000000000000000000: CC_MUX_REG_TO_BUS_OUT = REG_TO_MUX_R31;
		38'b00000100000000000000000000000000000000: CC_MUX_REG_TO_BUS_OUT = REG_TO_MUX_R32;
		38'b00001000000000000000000000000000000000: CC_MUX_REG_TO_BUS_OUT = REG_TO_MUX_R33;
		38'b00010000000000000000000000000000000000: CC_MUX_REG_TO_BUS_OUT = REG_TO_MUX_R34;
		38'b00100000000000000000000000000000000000: CC_MUX_REG_TO_BUS_OUT = REG_TO_MUX_R35;
		38'b01000000000000000000000000000000000000: CC_MUX_REG_TO_BUS_OUT = REG_TO_MUX_R36;
		38'b10000000000000000000000000000000000000: CC_MUX_REG_TO_BUS_OUT = REG_TO_MUX_R37;
		default : CC_MUX_REG_TO_BUS_OUT = 0;
		endcase
	end
endmodule
